`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:54:13 03/14/2014 
// Design Name: 
// Module Name:    ts_diff 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ts_diff(

clk,
rst,

ts_din,
ts_din_en,

ts_dout,
ts_dout_en



    );


input  			clk;
input			rst;
input	[32:0]	ts_din;
input 			ts_din_en;


output 	[32:0]	ts_dout;
output 			ts_dout_en;

reg 	[32:0]	ts_dout;
reg 			ts_dout_en;

reg 	[7:0]	ts_cnt;
reg 	[32:0]	ts_din_r1,ts_din_r2,ts_din_r3,ts_din_r4;
reg 			ts_din_en_r1,ts_din_en_r2;
reg 			send_flag;

always @(posedge clk)
begin
ts_din_en_r1<=ts_din_en;
ts_din_en_r2<=ts_din_en_r1;
ts_din_r1	<=ts_din;
ts_din_r2	<=ts_din_r1;
ts_din_r3	<=ts_din_r2;
ts_din_r4	<=ts_din_r3;
end

always@(posedge clk)
begin
if(rst)
	ts_cnt	<=0;
else if(ts_din_en | ts_din_en_r2)
	ts_cnt	<=ts_cnt+1;
else 
	ts_cnt	<=0;
end

always@(posedge clk)
begin
if(rst)
send_flag	<=0;
else if(ts_cnt==3 && ts_din[31:24]==8'h47)
	send_flag	<=1;
else if(ts_cnt	>1)
	send_flag	<=send_flag;
else 
send_flag	<=0;
end




always@(posedge clk)
begin
if(rst)
begin
ts_dout	<=0;
ts_dout_en	<=0;
end
else if(send_flag)
begin
ts_dout <=ts_din_r4;
ts_dout_en	<=1;
end
else 
begin
ts_dout	<=0;
ts_dout_en	<=0;
end
end

endmodule

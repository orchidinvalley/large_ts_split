`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:56:51 09/23/2019
// Design Name:   tsmf_split_v1
// Module Name:   E:/FPGA_pro/pcie_4gbe/tsmf_split_v1_test.v
// Project Name:  pcie_4g_gbe
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: tsmf_split_v1
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tsmf_split_v1_test;

	// Inputs
	reg clk;
	reg rst;
	reg [31:0] ts_din;
	reg ts_din_en;
	reg [7:0] freq_con_din;
	reg freq_con_din_en;
	reg [7:0] channel_din;
	reg channel_din_en;

	// Outputs
	wire ts_ram_wr;
	wire [511:0] ts_ram_wdata;
	wire test_flag;

	// Instantiate the Unit Under Test (UUT)
	tsmf_split_v1 uut (
		.clk(clk), 
		.rst(rst), 
		.ts_din(ts_din), 
		.ts_din_en(ts_din_en), 
		.freq_con_din(freq_con_din), 
		.freq_con_din_en(freq_con_din_en), 
		.channel_din(channel_din), 
		.channel_din_en(channel_din_en), 
		.ts_ram_wr(ts_ram_wr), 
		.ts_ram_wdata(ts_ram_wdata), 
		.test_flag(test_flag)
	);

	reg[31:0]i;

  reg[3:0]cnt=0;
  reg[31:0]rand;


	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 0;
		ts_din = 0;
		ts_din_en = 0;
		freq_con_din = 0;
		freq_con_din_en = 0;
		channel_din = 0;
		channel_din_en = 0;

		// Wait 100 ns for global reset to finish
		#1000;
        
    #2 rst =1;
		// Wait 100 ns for global reset to finish
		#1000;
		
			rst=0;
			
			
		
			
		#1000;
		
		#10 freq_con_din_en=1;
		freq_con_din=00;
		#10 freq_con_din=00;
		#10 freq_con_din=1;
		#10 freq_con_din=0;
		#10 freq_con_din=80;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;		
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din=0;
		#10 freq_con_din_en=0;
		
		
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
        #1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;    
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
			#1000;
		
		ts_send();
		cnt=cnt+1;
		#1000;
		
		ts_send();
		cnt=cnt+1;
		// Add stimulus here

	end
	
	always #5 clk=~clk;
	
	task ts_send();
	begin
	rand={$random}%16;
	#10 ts_din_en=1;
  ts_din=1;
  #10 ts_din={28'h4710010,cnt};
  
  for(i=1;i<47;i=i+1)
  #10 ts_din=i;
 	#10 ts_din_en=0;
 	ts_din=0;
 	
 	#100;
	end
	endtask
      
endmodule

